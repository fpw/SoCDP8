-- Part of SoCDP8, Copyright by Folke Will, 2019
-- Licensed under CERN Open Hardware Licence v1.2
-- See HW_LICENSE for details
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

use work.socdp8_package.all;
use work.pidp8_console_package.all;

entity pdp8 is
    generic (
        clk_frq: natural
    );
    port (
        clk: in std_logic;
        rst: in std_logic;
        
        -- Console connection
        leds: out pdp8i_leds;
        switches: in pdp8i_switches;

        -- to be connected to the external memory
        ext_mem_in: in ext_mem_in;
        ext_mem_out: out ext_mem_out
    );
end pdp8;

architecture Behavioral of pdp8 is
    -- whether to generate continuous memory cycles
    signal run: std_logic;

    -- current major state
    signal state: pdp8_state;

    -- interrupt on FF
    signal ion: std_logic;
    
    -- the manual preset signal clears the major state
    signal manual_preset: std_logic;
    -- the initialize signal clears several circuits
    signal initialize: std_logic;

    -- interconnect wires
    --- from manual timing generator
    signal mft: manual_function_time;
    signal mftp: std_logic;
    signal mfts0: std_logic;
    --- from memory
    signal strobe: std_logic;
    signal sense: std_logic_vector(11 downto 0);
    signal mem_start: std_logic;
    signal mem_done: std_logic;
    --- from register network
    signal carry_insert, no_shift, link: std_logic;
    signal pc, ma, mb, ac, mem: std_logic_vector(11 downto 0);
    signal inst: pdp8_instruction;
    signal ac_enable, pc_enable, ma_enable, mem_enable, sr_enable: std_logic;
    signal ac_load, pc_load, ma_load, mb_load: std_logic;
begin

manual_timing_inst: entity work.manual_timing
generic map (
    clk_frq => clk_frq
)
port map (
    clk => clk,
    rst => rst,
    run => run,
    
    key_load => switches.load,
    key_start => switches.start,
    key_ex => switches.exam,
    key_dep => switches.dep,
    key_cont => switches.cont,
    
    mfts0 => mfts0,
    mftp => mftp,
    mft => mft
);

regs: entity work.registers
port map (
    clk => clk,
    rst => rst,
    
    sr => switches.swr,
    sense => sense,
    
    initialize => initialize,
    carry_insert => carry_insert,
    no_shift => no_shift,
    
    pc_o => pc,
    ma_o => ma,
    mb_o => mb,
    ac_o => ac,
    link_o => link,
    inst_o => inst,
    
    ac_enable => ac_enable,
    pc_enable => pc_enable,
    ma_enable => ma_enable,
    mem_enable => mem_enable,
    sr_enable => sr_enable,
    
    ac_load => ac_load,
    pc_load => pc_load,
    ma_load => ma_load,
    mb_load => mb_load
);

mem_control: entity work.memory_control
generic map (
    clk_frq => clk_frq
)
port map (
    clk => clk,
    rst => rst,
    mem_addr => ma,
    field => "000",
    mem_start => mem_start,
    mem_done => mem_done,
    strobe => strobe,
    sense => sense,
    mem_buf => mb,
    ext_mem_in => ext_mem_in,
    ext_mem_out => ext_mem_out
);

time_states: process
begin
    wait until rising_edge(clk);
    
    -- reset pulse signals
    --- internal
    manual_preset <= '0';
    initialize <= '0';

    --- registers    
    no_shift <= '1';
    carry_insert <= '0';
    ac_enable <= '0';
    pc_enable <= '0';
    ma_enable <= '0';
    mem_enable <= '0';
    sr_enable <= '0';
    ac_load <= '0';
    pc_load <= '0';
    ma_load <= '0';
    mb_load <= '0';
    
    if mftp = '1' then
        case mft is
            when MFT_NONE =>
            when MFT1 =>
            when MFT2 =>
            when MFT3 =>
        end case;
    end if;
    
    -- generated by LA, START, EX, DEP
    if manual_preset = '1' then
        run <= '0';
        state <= STATE_MANUAL;
        ion <= '0';
    end if;

    -- generated by start switch
    if initialize = '1' then
        state <= STATE_FETCH;
        ion <= '0';
    end if;

    if rst = '1' then
        run <= '0';
        state <= STATE_MANUAL;
        ion <= '0';
    end if;
end process;

leds.pc <= pc;
leds.mem_addr <= ma;
leds.mem_buf <= mb;
leds.accu <= ac;
leds.link <= link;

leds.state <= state;
leds.instruction <= inst;
leds.ion <= ion;
leds.run <= run;

end Behavioral;
